//�ṹ��������ʽ����ģ�������Ϊ������ʽ��ʵ������4.1�Ĳ�һ�µ�·������Ϊ����ߵ�3���������أ����Ϊ����ߵ�LED�ơ�

`timescale 1ns / 1ps	

module not_gate(
    input a,
    output reg f                               
);
    always @(*)                        //��Ϊ������ʽ
    begin
        f <= ~a; 
    end
endmodule

module or_gate(
    input a,
    input b,
    output reg f                               
);
    always @(*)                        //��Ϊ������ʽ
    begin
        f <= a | b; 
    end
endmodule

module nand_gate(
    input a,
    input b,
    output reg f                               
);
    always @(*)                        //��Ϊ������ʽ
    begin
        f <= ~(a & b); 
    end
endmodule

module example_4_1(
    input sw_pin[7:0],                               		 //8����������
    output [15:0] led_pin    		 	//16��led��            
);
    wire p1, p2, p3, p4, p5;
    not_gate U1(.a(sw_pin[0]),.f(p1));				//�ṹ��������ʽ
    or_gate U2(.a(sw_pin[1]),.b(sw_pin[2]),.f(p2));			//�ṹ��������ʽ
    nand_gate U3(.a(sw_pin[1]),.b(sw_pin[2]),.f(p3));		//�ṹ��������ʽ
    nand_gate U4(.a(p1),.b(p2),.f(p4));				//�ṹ��������ʽ
    nand_gate U5(.a(p3),.b(sw_pin[0]),.f(p5));			//�ṹ��������ʽ
    nand_gate U6(.a(p4),.b(p5),.f(led_pin[0]));			//�ṹ��������ʽ
endmodule
//������Ϊ������ʽʵ���߶���ʾ������������AΪ����������ߵ�4���������أ�����BΪ���������ұߵ�4���������أ����Ϊ�������ϵ�8������ܣ����4����ӦA��ʮ������ֵ���ұ�4����ӦB��ʮ������ֵ����

`timescale 1ns / 1ps

module segment_display_decoder(
    input [7:0] sw_pin,					//8����������
    output [7:0] seg_data_0_pin, seg_data_1_pin, seg_cs_pin		//8�������
);

    reg [7:0] seg0, seg1;

    always @(*)                        //��Ϊ������ʽ
    begin
                case({sw_pin[0],sw_pin[1],sw_pin[2],sw_pin[3]})
	               0: 	seg0 <= 8'h3f;			    //  ��ߵ�4���������ʾ��0��
	               1: 	seg0 <= 8'h06;			    //  ��ߵ�4���������ʾ��1��
	               2: 	seg0 <= 8'h5b;			    //  ��ߵ�4���������ʾ��2��
	               3: 	seg0 <= 8'h4f;			    //  ��ߵ�4���������ʾ��3��
	               4: 	seg0 <= 8'h66;			    //  ��ߵ�4���������ʾ��4��
	               5: 	seg0 <= 8'h6d;			    //  ��ߵ�4���������ʾ��5��
	               6: 	seg0 <= 8'h7d;			    //  ��ߵ�4���������ʾ��6��
	               7: 	seg0 <= 8'h07;			    //  ��ߵ�4���������ʾ��7��
	               8: 	seg0 <= 8'h7f;			    //  ��ߵ�4���������ʾ��8��
	               9: 	seg0 <= 8'h6f;			    //  ��ߵ�4���������ʾ��9��
	               10: 	seg0 <= 8'h77;			    //  ��ߵ�4���������ʾ��A��
	               11: 	seg0 <= 8'h7c;			    //  ��ߵ�4���������ʾ��b��
	               12: 	seg0 <= 8'h39;			    //  ��ߵ�4���������ʾ��c��
	               13: 	seg0 <= 8'h5e;			    //  ��ߵ�4���������ʾ��d��
	               14: 	seg0 <= 8'h79;			    //  ��ߵ�4���������ʾ��E��
	               15: 	seg0 <= 8'h71;			    //  ��ߵ�4���������ʾ��F��
	               default:     seg0 <= 8'h00;			    //  ��ߵ�4�������ȫ��
                endcase

                case({sw_pin[4],sw_pin[5],sw_pin[6],sw_pin[7]})
	               0: 	seg1 <= 8'h3f;			    //  �ұߵ�4���������ʾ��0��
	               1: 	seg1 <= 8'h06;			    //  �ұߵ�4���������ʾ��1��
	               2: 	seg1 <= 8'h5b;			    //  �ұߵ�4���������ʾ��2��
	               3: 	seg1 <= 8'h4f;			    //  �ұߵ�4���������ʾ��3��
	               4: 	seg1 <= 8'h66;			    //  �ұߵ�4���������ʾ��4��
	               5: 	seg1 <= 8'h6d;			    //  �ұߵ�4���������ʾ��5��
	               6: 	seg1 <= 8'h7d;			    //  �ұߵ�4���������ʾ��6��
	               7: 	seg1 <= 8'h07;			    //  �ұߵ�4���������ʾ��7��
	               8: 	seg1 <= 8'h7f;			    //  �ұߵ�4���������ʾ��8��
	               9: 	seg1 <= 8'h6f;			    //  �ұߵ�4���������ʾ��9��
	               10: 	seg1 <= 8'h77;			    //  �ұߵ�4���������ʾ��A��
	               11: 	seg1 <= 8'h7c;			    //  �ұߵ�4���������ʾ��b��
	               12: 	seg1 <= 8'h39;			    //  �ұߵ�4���������ʾ��c��
	               13: 	seg1 <= 8'h5e;			    //  �ұߵ�4���������ʾ��d��
	               14: 	seg1 <= 8'h79;			    //  �ұߵ�4���������ʾ��E��
	               15: 	seg1 <= 8'h71;			    //  �ұߵ�4���������ʾ��F��
	               default:     seg1 <= 8'h00;			    //  ��ߵ�4�������ȫ��
                endcase
    end

    assign seg_data_0_pin = seg0;		//���4������ܵ�8����
    assign seg_data_1_pin = seg1;		//�ұ�4������ܵ�8����
    assign seg_cs_pin = 8'hff;                              	//8������ܵ�8��λ

endmodule